
-- This component is a decimal counter based on the input I as regard to an internal time reference

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CPT_decimal is
  Port ( CLK : in  STD_LOGIC;
         RAZ : in  STD_LOGIC;
         I : in STD_LOGIC;
         Q: out INTEGER);
end CPT_decimal;

architecture Behavioral of CPT_decimal is
signal internalQ : INTEGER := 0; -- internal signal of output Q
signal internalCLK : STD_LOGIC; -- Internal clock, generated by the clock manager
							    -- This is the time reference to count

component clock_manager -- Declaration of the clock manager
    Port ( MAINCLK : in STD_LOGIC;
           BAUDRATE : in INTEGER;
           CLKOUT : out STD_LOGIC);
end component;

begin
Q <= internalQ;

-- Clock generator
CLKMGT : clock_manager port map (CLK, 1000000, internalCLK);
-- We will take baudrate=1000000 for the test bench (for faster simulation calcul)
-- and baudrate=2 to test on ZBoard (2 evaluations per second)

process (I, RAZ, internalCLK)
begin
if RAZ='1' then internalQ <= 0;
elsif (internalCLK'event and internalCLK='1') then
	if I='1' then
		if internalQ=9999 then internalQ <= 0;
		else internalQ <= (internalQ+1);
		end if;
    end if;
   end if;
end process;
end Behavioral;
